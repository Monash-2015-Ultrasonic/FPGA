module hex_output(
	input 	[15:0]	data,
	output 	[8:0] 	display
	);
	
	
	
	
	
endmodule
