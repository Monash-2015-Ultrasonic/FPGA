// test_qsys.v

// Generated using ACDS version 13.0sp1 232 at 2015.03.22.20:48:01

`timescale 1 ps / 1 ps
module test_qsys (
		input  wire  clk_qsys_50_clk,     //    clk_qsys_50.clk
		input  wire  reset_reset_n,       //          reset.reset_n
		input  wire  spi_0_external_MISO, // spi_0_external.MISO
		output wire  spi_0_external_MOSI, //               .MOSI
		output wire  spi_0_external_SCLK, //               .SCLK
		input wire  spi_0_external_SS_n  //               .SS_n
	);

	wire    rst_controller_reset_out_reset; // rst_controller:reset_out -> spi_0:reset_n

	test_qsys_spi_0 spi_0 (
		.clk           (clk_qsys_50_clk),                 //              clk.clk
		.reset_n       (~rst_controller_reset_out_reset), //            reset.reset_n
		.data_from_cpu (),                                // spi_control_port.writedata
		.data_to_cpu   (),                                //                 .readdata
		.mem_addr      (),                                //                 .address
		.read_n        (),                                //                 .read_n
		.spi_select    (spi_0_external_SS_n),                                //                 .chipselect
		.write_n       (),                                //                 .write_n
		.irq           (),                                //              irq.irq
		.MISO          (spi_0_external_MISO),             //         external.export
		.MOSI          (spi_0_external_MOSI),             //                 .export
		.SCLK          (spi_0_external_SCLK),             //                 .export
		.SS_n          ()              //                 .export
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                 // reset_in0.reset
		.clk        (clk_qsys_50_clk),                //       clk.clk
		.reset_out  (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req  (),                               // (terminated)
		.reset_in1  (1'b0),                           // (terminated)
		.reset_in2  (1'b0),                           // (terminated)
		.reset_in3  (1'b0),                           // (terminated)
		.reset_in4  (1'b0),                           // (terminated)
		.reset_in5  (1'b0),                           // (terminated)
		.reset_in6  (1'b0),                           // (terminated)
		.reset_in7  (1'b0),                           // (terminated)
		.reset_in8  (1'b0),                           // (terminated)
		.reset_in9  (1'b0),                           // (terminated)
		.reset_in10 (1'b0),                           // (terminated)
		.reset_in11 (1'b0),                           // (terminated)
		.reset_in12 (1'b0),                           // (terminated)
		.reset_in13 (1'b0),                           // (terminated)
		.reset_in14 (1'b0),                           // (terminated)
		.reset_in15 (1'b0)                            // (terminated)
	);

endmodule
