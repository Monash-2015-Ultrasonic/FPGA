module inSumSquare(
	input SYS_CLK,
	input [11:0] inValue,
	input validCondition,
	output reg [23:0] outValue
	);

reg [11:0] x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200, x201, x202, x203, x204, x205, x206, x207, x208, x209, x210, x211, x212, x213, x214, x215, x216, x217, x218, x219, x220, x221, x222, x223, x224, x225, x226, x227, x228, x229, x230, x231, x232, x233, x234, x235, x236, x237, x238, x239, x240, x241, x242, x243, x244, x245, x246, x247, x248, x249, x250, x251, x252, x253, x254, x255, x256, x257, x258, x259;


always @(posedge SYS_CLK) begin
	if (validCondition) begin
		x0 <= inValue;
		x1 <= x0;
		x2 <= x1;
		x3 <= x2;
		x4 <= x3;
		x5 <= x4;
		x6 <= x5;
		x7 <= x6;
		x8 <= x7;
		x9 <= x8;
		x10 <= x9;
		x11 <= x10;
		x12 <= x11;
		x13 <= x12;
		x14 <= x13;
		x15 <= x14;
		x16 <= x15;
		x17 <= x16;
		x18 <= x17;
		x19 <= x18;
		x20 <= x19;
		x21 <= x20;
		x22 <= x21;
		x23 <= x22;
		x24 <= x23;
		x25 <= x24;
		x26 <= x25;
		x27 <= x26;
		x28 <= x27;
		x29 <= x28;
		x30 <= x29;
		x31 <= x30;
		x32 <= x31;
		x33 <= x32;
		x34 <= x33;
		x35 <= x34;
		x36 <= x35;
		x37 <= x36;
		x38 <= x37;
		x39 <= x38;
		x40 <= x39;
		x41 <= x40;
		x42 <= x41;
		x43 <= x42;
		x44 <= x43;
		x45 <= x44;
		x46 <= x45;
		x47 <= x46;
		x48 <= x47;
		x49 <= x48;
		x50 <= x49;
		x51 <= x50;
		x52 <= x51;
		x53 <= x52;
		x54 <= x53;
		x55 <= x54;
		x56 <= x55;
		x57 <= x56;
		x58 <= x57;
		x59 <= x58;
		x60 <= x59;
		x61 <= x60;
		x62 <= x61;
		x63 <= x62;
		x64 <= x63;
		x65 <= x64;
		x66 <= x65;
		x67 <= x66;
		x68 <= x67;
		x69 <= x68;
		x70 <= x69;
		x71 <= x70;
		x72 <= x71;
		x73 <= x72;
		x74 <= x73;
		x75 <= x74;
		x76 <= x75;
		x77 <= x76;
		x78 <= x77;
		x79 <= x78;
		x80 <= x79;
		x81 <= x80;
		x82 <= x81;
		x83 <= x82;
		x84 <= x83;
		x85 <= x84;
		x86 <= x85;
		x87 <= x86;
		x88 <= x87;
		x89 <= x88;
		x90 <= x89;
		x91 <= x90;
		x92 <= x91;
		x93 <= x92;
		x94 <= x93;
		x95 <= x94;
		x96 <= x95;
		x97 <= x96;
		x98 <= x97;
		x99 <= x98;
		x100 <= x99;
		x101 <= x100;
		x102 <= x101;
		x103 <= x102;
		x104 <= x103;
		x105 <= x104;
		x106 <= x105;
		x107 <= x106;
		x108 <= x107;
		x109 <= x108;
		x110 <= x109;
		x111 <= x110;
		x112 <= x111;
		x113 <= x112;
		x114 <= x113;
		x115 <= x114;
		x116 <= x115;
		x117 <= x116;
		x118 <= x117;
		x119 <= x118;
		x120 <= x119;
		x121 <= x120;
		x122 <= x121;
		x123 <= x122;
		x124 <= x123;
		x125 <= x124;
		x126 <= x125;
		x127 <= x126;
		x128 <= x127;
		x129 <= x128;
		x130 <= x129;
		x131 <= x130;
		x132 <= x131;
		x133 <= x132;
		x134 <= x133;
		x135 <= x134;
		x136 <= x135;
		x137 <= x136;
		x138 <= x137;
		x139 <= x138;
		x140 <= x139;
		x141 <= x140;
		x142 <= x141;
		x143 <= x142;
		x144 <= x143;
		x145 <= x144;
		x146 <= x145;
		x147 <= x146;
		x148 <= x147;
		x149 <= x148;
		x150 <= x149;
		x151 <= x150;
		x152 <= x151;
		x153 <= x152;
		x154 <= x153;
		x155 <= x154;
		x156 <= x155;
		x157 <= x156;
		x158 <= x157;
		x159 <= x158;
		x160 <= x159;
		x161 <= x160;
		x162 <= x161;
		x163 <= x162;
		x164 <= x163;
		x165 <= x164;
		x166 <= x165;
		x167 <= x166;
		x168 <= x167;
		x169 <= x168;
		x170 <= x169;
		x171 <= x170;
		x172 <= x171;
		x173 <= x172;
		x174 <= x173;
		x175 <= x174;
		x176 <= x175;
		x177 <= x176;
		x178 <= x177;
		x179 <= x178;
		x180 <= x179;
		x181 <= x180;
		x182 <= x181;
		x183 <= x182;
		x184 <= x183;
		x185 <= x184;
		x186 <= x185;
		x187 <= x186;
		x188 <= x187;
		x189 <= x188;
		x190 <= x189;
		x191 <= x190;
		x192 <= x191;
		x193 <= x192;
		x194 <= x193;
		x195 <= x194;
		x196 <= x195;
		x197 <= x196;
		x198 <= x197;
		x199 <= x198;
		x200 <= x199;
		x201 <= x200;
		x202 <= x201;
		x203 <= x202;
		x204 <= x203;
		x205 <= x204;
		x206 <= x205;
		x207 <= x206;
		x208 <= x207;
		x209 <= x208;
		x210 <= x209;
		x211 <= x210;
		x212 <= x211;
		x213 <= x212;
		x214 <= x213;
		x215 <= x214;
		x216 <= x215;
		x217 <= x216;
		x218 <= x217;
		x219 <= x218;
		x220 <= x219;
		x221 <= x220;
		x222 <= x221;
		x223 <= x222;
		x224 <= x223;
		x225 <= x224;
		x226 <= x225;
		x227 <= x226;
		x228 <= x227;
		x229 <= x228;
		x230 <= x229;
		x231 <= x230;
		x232 <= x231;
		x233 <= x232;
		x234 <= x233;
		x235 <= x234;
		x236 <= x235;
		x237 <= x236;
		x238 <= x237;
		x239 <= x238;
		x240 <= x239;
		x241 <= x240;
		x242 <= x241;
		x243 <= x242;
		x244 <= x243;
		x245 <= x244;
		x246 <= x245;
		x247 <= x246;
		x248 <= x247;
		x249 <= x248;
		x250 <= x249;
		x251 <= x250;
		x252 <= x251;
		x253 <= x252;
		x254 <= x253;
		x255 <= x254;
		x256 <= x255;
		x257 <= x256;
		x258 <= x257;
		x259 <= x258;
	end
end

always @(posedge SYS_CLK) begin
	if (validCondition) begin
		outValue <= x0*x0 + x1*x1 + x2*x2 + x3*x3 + x4*x4 + x5*x5 + x6*x6 + x7*x7 + x8*x8 + x9*x9 + x10*x10 + x11*x11 + x12*x12 + x13*x13 + x14*x14 + x15*x15 + x16*x16 + x17*x17 + x18*x18 + x19*x19 + x20*x20 + x21*x21 + x22*x22 + x23*x23 + x24*x24 + x25*x25 + x26*x26 + x27*x27 + x28*x28 + x29*x29 + x30*x30 + x31*x31 + x32*x32 + x33*x33 + x34*x34 + x35*x35 + x36*x36 + x37*x37 + x38*x38 + x39*x39 + x40*x40 + x41*x41 + x42*x42 + x43*x43 + x44*x44 + x45*x45 + x46*x46 + x47*x47 + x48*x48 + x49*x49 + x50*x50 + x51*x51 + x52*x52 + x53*x53 + x54*x54 + x55*x55 + x56*x56 + x57*x57 + x58*x58 + x59*x59 + x60*x60 + x61*x61 + x62*x62 + x63*x63 + x64*x64 + x65*x65 + x66*x66 + x67*x67 + x68*x68 + x69*x69 + x70*x70 + x71*x71 + x72*x72 + x73*x73 + x74*x74 + x75*x75 + x76*x76 + x77*x77 + x78*x78 + x79*x79 + x80*x80 + x81*x81 + x82*x82 + x83*x83 + x84*x84 + x85*x85 + x86*x86 + x87*x87 + x88*x88 + x89*x89 + x90*x90 + x91*x91 + x92*x92 + x93*x93 + x94*x94 + x95*x95 + x96*x96 + x97*x97 + x98*x98 + x99*x99 + x100*x100 + x101*x101 + x102*x102 + x103*x103 + x104*x104 + x105*x105 + x106*x106 + x107*x107 + x108*x108 + x109*x109 + x110*x110 + x111*x111 + x112*x112 + x113*x113 + x114*x114 + x115*x115 + x116*x116 + x117*x117 + x118*x118 + x119*x119 + x120*x120 + x121*x121 + x122*x122 + x123*x123 + x124*x124 + x125*x125 + x126*x126 + x127*x127 + x128*x128 + x129*x129 + x130*x130 + x131*x131 + x132*x132 + x133*x133 + x134*x134 + x135*x135 + x136*x136 + x137*x137 + x138*x138 + x139*x139 + x140*x140 + x141*x141 + x142*x142 + x143*x143 + x144*x144 + x145*x145 + x146*x146 + x147*x147 + x148*x148 + x149*x149 + x150*x150 + x151*x151 + x152*x152 + x153*x153 + x154*x154 + x155*x155 + x156*x156 + x157*x157 + x158*x158 + x159*x159 + x160*x160 + x161*x161 + x162*x162 + x163*x163 + x164*x164 + x165*x165 + x166*x166 + x167*x167 + x168*x168 + x169*x169 + x170*x170 + x171*x171 + x172*x172 + x173*x173 + x174*x174 + x175*x175 + x176*x176 + x177*x177 + x178*x178 + x179*x179 + x180*x180 + x181*x181 + x182*x182 + x183*x183 + x184*x184 + x185*x185 + x186*x186 + x187*x187 + x188*x188 + x189*x189 + x190*x190 + x191*x191 + x192*x192 + x193*x193 + x194*x194 + x195*x195 + x196*x196 + x197*x197 + x198*x198 + x199*x199 + x200*x200 + x201*x201 + x202*x202 + x203*x203 + x204*x204 + x205*x205 + x206*x206 + x207*x207 + x208*x208 + x209*x209 + x210*x210 + x211*x211 + x212*x212 + x213*x213 + x214*x214 + x215*x215 + x216*x216 + x217*x217 + x218*x218 + x219*x219 + x220*x220 + x221*x221 + x222*x222 + x223*x223 + x224*x224 + x225*x225 + x226*x226 + x227*x227 + x228*x228 + x229*x229 + x230*x230 + x231*x231 + x232*x232 + x233*x233 + x234*x234 + x235*x235 + x236*x236 + x237*x237 + x238*x238 + x239*x239 + x240*x240 + x241*x241 + x242*x242 + x243*x243 + x244*x244 + x245*x245 + x246*x246 + x247*x247 + x248*x248 + x249*x249 + x250*x250 + x251*x251 + x252*x252 + x253*x253 + x254*x254 + x255*x255 + x256*x256 + x257*x257 + x258*x258 + x259*x259;
	end
	else begin
		outValue <= outValue;
	end
end

endmodule
