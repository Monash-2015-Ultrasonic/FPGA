module SignalGen(
	
	
	);
	
	
	
	//
	// High
	// Wait 12.5us
	// Low
	// x4
	
	
endmodule	
